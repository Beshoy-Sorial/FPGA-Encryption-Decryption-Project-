module InvShiftRows(input [0:127]state,output  [0:127]out);

assign out[0:127] = { state[0:7] , state[104:111] ,state[80:87] , state[56:63] 
                    , state[32:39] , state[8:15] , state[112:119] , state[88:95]  
                    , state[64:71] , state[40:47] , state[16:23] , state[120:127] 
                    , state[96:103] , state[72:79] , state[48:55] , state[24:31]  } ; 


endmodule

