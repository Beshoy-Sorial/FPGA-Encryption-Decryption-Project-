module Manager(input s1,s2,reset,clk,output reg L1,L2,L3,output [6:0]H,T,O);

integer i = 0;
wire [127:0] out1;
wire [127:0] out2;
wire [127:0] out3;
wire [127:0] out4;
wire [127:0] out5;
wire [127:0] out6;
reg  [127:0] final;	//Final Output ================> Put last 8 bits [7:0] in BCD #(BCD wihtout clk)
wire [11:0] bcd;


bin2bcd b(final [7:0],bcd);

segment7 s5(bcd[11:8],H);
segment7 s6(bcd[7:4],T);
segment7 s7(bcd[3:0],O);

wire [127:0] in = 128'h_00112233445566778899aabbccddeeff;					

wire [127:0] k1 = 128'h_000102030405060708090a0b0c0d0e0f;					
wire [191:0] k2 = 192'h_000102030405060708090a0b0c0d0e0f1011121314151617;			
wire [255:0] k3 = 256'h_000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f ;	 

  Encrypt #(4,10) E1 (clk,reset,in,k1,out1);
  Encrypt #(6,12) E2 (clk,reset,in,k2,out2);
  Encrypt #(8,14) E3 (clk,reset,in,k3,out3);
  Decrypt #(4,10) D1 (out1,k1,out4,clk,reset);
  Decrypt #(6,12) D2 (out2,k2,out5,clk,reset);
  Decrypt #(8,14) D3 (out3,k3,out6,clk,reset);

always @(posedge clk or posedge reset) begin
if (reset) i = 0;
else i = i + 1;
end


always @(*) begin

if (!s1 && !s2) begin 

if (i <= 11)
final <= out1; 
else
final <= out4;
end
else if (s1 && !s2) begin 

if (i <= 13)
final <= out2; 
else
final <= out5;
end
else if (!s1 && s2) begin 

if (i <= 15)
final <= out3; 
else
final <= out6;
end



if( out4== in) begin
L1<=1;
end
else begin
L1<=0;
end

if( out5== in) begin
L2<=1;
end
else begin
L2<=0;
end

if(out6 == in) begin
L3<=1;
end
else begin
L3<=0;
end




end

 
endmodule